
module this_clock (
	oscena,
	clkout);	

	input		oscena;
	output		clkout;
endmodule
