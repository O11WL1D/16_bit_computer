-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Thu May 18 16:17:16 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY control_mod IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        general : IN STD_LOGIC := '0';
        ram_write_enable : OUT STD_LOGIC;
        progcountTOram : OUT STD_LOGIC;
        programcontincrement : OUT STD_LOGIC;
        programcontenable : OUT STD_LOGIC;
        state0 : OUT STD_LOGIC;
        state1 : OUT STD_LOGIC;
        state2 : OUT STD_LOGIC;
        super0 : OUT STD_LOGIC;
        super1 : OUT STD_LOGIC
    );
END control_mod;

ARCHITECTURE BEHAVIOR OF control_mod IS
    TYPE type_fstate IS (i1m0,i1m1,wait0,i2m0resetpc,i3m0readram,state4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,general)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= wait0;
            ram_write_enable <= '0';
            progcountTOram <= '0';
            programcontincrement <= '0';
            programcontenable <= '0';
            state0 <= '0';
            state1 <= '0';
            state2 <= '0';
            super0 <= '0';
            super1 <= '0';
        ELSE
            ram_write_enable <= '0';
            progcountTOram <= '0';
            programcontincrement <= '0';
            programcontenable <= '0';
            state0 <= '0';
            state1 <= '0';
            state2 <= '0';
            super0 <= '0';
            super1 <= '0';
            CASE fstate IS
                WHEN i1m0 =>
                    IF ((general = '1')) THEN
                        reg_fstate <= i1m1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= i1m0;
                    END IF;

                    ram_write_enable <= '0';

                    programcontenable <= '1';

                    state0 <= '1';

                    programcontincrement <= '1';

                    state2 <= '0';

                    super1 <= '0';

                    super0 <= '1';

                    progcountTOram <= '0';

                    state1 <= '0';
                WHEN i1m1 =>
                    IF ((general = '1')) THEN
                        reg_fstate <= wait0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= i1m1;
                    END IF;

                    ram_write_enable <= '1';

                    state0 <= '0';

                    state2 <= '0';

                    super1 <= '0';

                    super0 <= '1';

                    progcountTOram <= '1';

                    state1 <= '1';
                WHEN wait0 =>
                    IF ((general = '1')) THEN
                        reg_fstate <= i1m0;
                    ELSIF ((general = '0')) THEN
                        reg_fstate <= i2m0resetpc;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= wait0;
                    END IF;

                    ram_write_enable <= '0';

                    state0 <= '0';

                    state2 <= '0';

                    super1 <= '0';

                    super0 <= '0';

                    state1 <= '0';
                WHEN i2m0resetpc =>
                    IF ((general = '0')) THEN
                        reg_fstate <= i3m0readram;
                    ELSIF ((general = '1')) THEN
                        reg_fstate <= wait0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= i2m0resetpc;
                    END IF;

                    ram_write_enable <= '0';

                    programcontenable <= '0';

                    state0 <= '0';

                    programcontincrement <= '1';

                    state2 <= '0';

                    super1 <= '1';

                    super0 <= '0';

                    progcountTOram <= '0';

                    state1 <= '0';
                WHEN i3m0readram =>
                    IF ((general = '0')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= i3m0readram;
                    END IF;

                    ram_write_enable <= '0';

                    programcontenable <= '0';
                    programcontenable <= '0';

                    state0 <= '0';

                    programcontincrement <= '0';

                    progcountTOram <= '1';
                WHEN state4 =>
                    IF ((general = '0')) THEN
                        reg_fstate <= i3m0readram;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    ram_write_enable <= '0';

                    programcontenable <= '1';

                    programcontincrement <= '1';

                    progcountTOram <= '0';
                WHEN OTHERS => 
                    ram_write_enable <= 'X';
                    progcountTOram <= 'X';
                    programcontincrement <= 'X';
                    programcontenable <= 'X';
                    state0 <= 'X';
                    state1 <= 'X';
                    state2 <= 'X';
                    super0 <= 'X';
                    super1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
