-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.


-- Generated by Quartus Prime Version 20.1 (Build Build 720 11/11/2020)
-- Created on Thu May 18 16:01:21 2023

control_mod control_mod_inst
(
	.reset(reset_sig) ,	// input  reset_sig
	.clock(clock_sig) ,	// input  clock_sig
	.ram_write_enable(ram_write_enable_sig) ,	// output  ram_write_enable_sig
	.progcountTOram(progcountTOram_sig) ,	// output  progcountTOram_sig
	.programcontincrement(programcontincrement_sig) ,	// output  programcontincrement_sig
	.programcontenable(programcontenable_sig) ,	// output  programcontenable_sig
	.state0(state0_sig) ,	// output  state0_sig
	.state1(state1_sig) ,	// output  state1_sig
	.state2(state2_sig) ,	// output  state2_sig
	.super0(super0_sig) ,	// output  super0_sig
	.super1(super1_sig) 	// output  super1_sig
);

