LIBRARY ieee;
USE ieee.std_logic_1164.all ;




Entity bus_split_64 is

port(


b : in std_logic_vector(63 downto 0) ;



A0, 
A1, 
A2, 
A3, 
A4, 
A5, 
A6, 
A7, 
A8, 
A9, 
A10, 
A11, 
A12, 
A13, 
A14, 
A15, 
A16, 
A17, 
A18, 
A19, 
A20, 
A21, 
A22, 
A23, 
A24, 
A25, 
A26, 
A27, 
A28, 
A29, 
A30, 
A31, 
A32, 
A33, 
A34, 
A35, 
A36, 
A37, 
A38, 
A39, 
A40, 
A41, 
A42, 
A43, 
A44, 
A45, 
A46, 
A47, 
A48, 
A49, 
A50, 
A51, 
A52, 
A53, 
A54, 
A55, 
A56, 
A57, 
A58, 
A59, 
A60, 
A61, 
A62, 
A63 :out std_logic




 



-- last item cannot have a semicolon 



);


end bus_split_64 ;




ARCHITECTURE LogicFunc of bus_split_64 is
Begin 


A0<=	b(0); 
A1<=	b(1); 
A2<=	b(2); 
A3<=	b(3); 
A4<=	b(4); 
A5<=	b(5); 
A6<=	b(6); 
A7<=	b(7); 
A8<=	b(8); 
A9<=	b(9); 
A10<=	b(10); 
A11<=	b(11); 
A12<=	b(12); 
A13<=	b(13); 
A14<=	b(14); 
A15<=	b(15); 
A16<=	b(16); 
A17<=	b(17); 
A18<=	b(18); 
A19<=	b(19); 
A20<=	b(20); 
A21<=	b(21); 
A22<=	b(22); 
A23<=	b(23); 
A24<=	b(24); 
A25<=	b(25); 
A26<=	b(26); 
A27<=	b(27); 
A28<=	b(28); 
A29<=	b(29); 
A30<=	b(30); 
A31<=	b(31); 
A32<=	b(32); 
A33<=	b(33); 
A34<=	b(34); 
A35<=	b(35); 
A36<=	b(36); 
A37<=	b(37); 
A38<=	b(38); 
A39<=	b(39); 
A40<=	b(40); 
A41<=	b(41); 
A42<=	b(42); 
A43<=	b(43); 
A44<=	b(44); 
A45<=	b(45); 
A46<=	b(46); 
A47<=	b(47); 
A48<=	b(48); 
A49<=	b(49); 
A50<=	b(50); 
A51<=	b(51); 
A52<=	b(52); 
A53<=	b(53); 
A54<=	b(54); 
A55<=	b(55); 
A56<=	b(56); 
A57<=	b(57); 
A58<=	b(58); 
A59<=	b(59); 
A60<=	b(60); 
A61<=	b(61); 
A62<=	b(62); 
A63<=	b(63); 








END LogicFunc ; 