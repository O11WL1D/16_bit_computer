-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Mon May 22 16:49:22 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY control_mod IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        test0 : IN STD_LOGIC := '0';
        test1 : IN STD_LOGIC := '0';
        ram_write_enable : OUT STD_LOGIC;
        progcountTOram : OUT STD_LOGIC;
        programcontincrement : OUT STD_LOGIC;
        programcontenable : OUT STD_LOGIC;
        saveRamAddr : OUT STD_LOGIC
    );
END control_mod;

ARCHITECTURE BEHAVIOR OF control_mod IS
    TYPE type_fstate IS (ramwrite0,ramwrite1,wait0,resetpc0,readram0,readram1);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,test0,test1)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= wait0;
            ram_write_enable <= '0';
            progcountTOram <= '0';
            programcontincrement <= '0';
            programcontenable <= '0';
            saveRamAddr <= '0';
        ELSE
            ram_write_enable <= '0';
            progcountTOram <= '0';
            programcontincrement <= '0';
            programcontenable <= '0';
            saveRamAddr <= '0';
            CASE fstate IS
                WHEN ramwrite0 =>
                    IF (((test0 = '1') AND NOT((test1 = '1')))) THEN
                        reg_fstate <= ramwrite1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ramwrite0;
                    END IF;

                    programcontincrement <= '1';

                    programcontenable <= '1';

                    progcountTOram <= '0';

                    ram_write_enable <= '0';
                WHEN ramwrite1 =>
                    IF (((test0 = '1') AND NOT((test1 = '1')))) THEN
                        reg_fstate <= wait0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ramwrite1;
                    END IF;

                    saveRamAddr <= '1';

                    progcountTOram <= '1';

                    ram_write_enable <= '1';
                WHEN wait0 =>
                    IF (((test0 = '1') AND NOT((test1 = '1')))) THEN
                        reg_fstate <= ramwrite0;
                    ELSIF ((NOT((test0 = '1')) AND (test1 = '1'))) THEN
                        reg_fstate <= resetpc0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= wait0;
                    END IF;

                    ram_write_enable <= '0';
                WHEN resetpc0 =>
                    IF ((NOT((test0 = '1')) AND (test1 = '1'))) THEN
                        reg_fstate <= readram0;
                    ELSIF (((test0 = '1') AND NOT((test1 = '1')))) THEN
                        reg_fstate <= wait0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= resetpc0;
                    END IF;

                    programcontincrement <= '1';

                    programcontenable <= '0';

                    progcountTOram <= '0';

                    ram_write_enable <= '0';
                WHEN readram0 =>
                    IF ((NOT((test0 = '1')) AND (test1 = '1'))) THEN
                        reg_fstate <= readram1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= readram0;
                    END IF;

                    programcontincrement <= '0';

                    saveRamAddr <= '1';

                    programcontenable <= '0';
                    programcontenable <= '0';

                    progcountTOram <= '1';

                    ram_write_enable <= '0';
                WHEN readram1 =>
                    IF ((NOT((test0 = '1')) AND (test1 = '1'))) THEN
                        reg_fstate <= readram0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= readram1;
                    END IF;

                    programcontincrement <= '1';

                    programcontenable <= '1';

                    progcountTOram <= '0';

                    ram_write_enable <= '0';
                WHEN OTHERS => 
                    ram_write_enable <= 'X';
                    progcountTOram <= 'X';
                    programcontincrement <= 'X';
                    programcontenable <= 'X';
                    saveRamAddr <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
