LIBRARY ieee ;
USE ieee.std_logic_1164.all ;




--let this be a lesson ; entity names cannot begin with a number :(





ENTITY  b16_en IS

PORT(

a : IN std_Logic_Vector(15 downto 0) ;

en : IN std_logic ;

f : OUT std_logic_VEctor(15 downto 0) 



-- last port should not contain a semicolon. :)

) ;

END b16_en; 









ARCHITECTURE LogicFunc of b16_en is

BEGIN 

f(     0    ) <= (a(   0     ) AND en) ;
f(     1    ) <= (a(   1     ) AND en) ;
f(     2    ) <= (a(   2     ) AND en) ;
f(     3    ) <= (a(   3     ) AND en) ;
f(     4    ) <= (a(   4     ) AND en) ;
f(     5    ) <= (a(   5     ) AND en) ;
f(     6    ) <= (a(   6     ) AND en) ;
f(     7    ) <= (a(   7     ) AND en) ;
f(     8    ) <= (a(   8     ) AND en) ;
f(     9    ) <= (a(   9     ) AND en) ;
f(10) <= (a(10) AND en) ;
f(11) <= (a(11) AND en) ;
f(12) <= (a(12) AND en) ;
f(13) <= (a(13) AND en) ;
f(14) <= (a(14) AND en) ;
f(15) <= (a(15) AND en) ;






end LogicFunc;
