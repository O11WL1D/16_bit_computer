
module testclock (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
