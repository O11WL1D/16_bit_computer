LIBRARY ieee;
USE ieee.std_logic_1164.all ;




Entity bus_split_32 is

port(


b : in std_logic_vector(31 downto 0) ;




A0, 
A1, 
A2, 
A3, 
A4, 
A5, 
A6, 
A7, 
A8, 
A9, 
A10, 
A11, 
A12, 
A13, 
A14, 
A15, 
A16, 
A17, 
A18, 
A19, 
A20, 
A21, 
A22, 
A23, 
A24, 
A25, 
A26, 
A27, 
A28, 
A29, 
A30, 
A31 :out std_logic




 



-- last item cannot have a semicolon 



);


end bus_split_32 ;




ARCHITECTURE LogicFunc of bus_split_32 is
Begin 


A0<=	b(0); 
A1<=	b(1); 
A2<=	b(2); 
A3<=	b(3); 
A4<=	b(4); 
A5<=	b(5); 
A6<=	b(6); 
A7<=	b(7); 
A8<=	b(8); 
A9<=	b(9); 
A10<=	b(10); 
A11<=	b(11); 
A12<=	b(12); 
A13<=	b(13); 
A14<=	b(14); 
A15<=	b(15); 
A16<=	b(16); 
A17<=	b(17); 
A18<=	b(18); 
A19<=	b(19); 
A20<=	b(20); 
A21<=	b(21); 
A22<=	b(22); 
A23<=	b(23); 
A24<=	b(24); 
A25<=	b(25); 
A26<=	b(26); 
A27<=	b(27); 
A28<=	b(28); 
A29<=	b(29); 
A30<=	b(30); 
A31<=	b(31); 









END LogicFunc ; 